library verilog;
use verilog.vl_types.all;
entity B is
    port(
        A_First         : in     vl_logic;
        A_Zero          : in     vl_logic;
        Zero            : in     vl_logic;
        BFlag           : out    vl_logic;
        instr           : in     vl_logic_vector(31 downto 26);
        addr            : in     vl_logic_vector(4 downto 0)
    );
end B;
