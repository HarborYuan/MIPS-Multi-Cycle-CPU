library verilog;
use verilog.vl_types.all;
entity PCUnit is
    port(
        \in\            : in     vl_logic_vector(31 downto 0);
        PC              : out    vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        sig             : in     vl_logic
    );
end PCUnit;
